module DataMemoryRegister(reset, clk);

input wire reset, clk;	




endmodule
