module DataMemoryRegister(reset, clk);

endmodule
