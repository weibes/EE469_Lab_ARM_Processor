module executeRegister(writeData, reset, clk);

endmodule
