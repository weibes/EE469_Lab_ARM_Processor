module registerFetchRegister(Data1, Data2, reset, clk);


endmodule
