module writebackRegister();


endmodule
